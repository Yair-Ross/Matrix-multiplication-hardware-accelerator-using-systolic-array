//
// Verilog Module Multiplexer_Accelarator_lib.memory_decoder
//
// Created:
//          by - rossy.UNKNOWN (SHOHAM)
//          at - 22:16:17 01/21/2024
//
// using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
//

`resetall
`timescale 1ns/10ps
module memory(clk_i, rst_ni, sp_mat_i, addr_i, read_i, write_i, wdata_i, flags_adder_i, flags_systolic_i, write_flag_i,strb_i, rdata_o, mod_o, 
 sp_read_o, sp_read_target_o, operand_A_o, operand_B_o, start_FMEM_o, write_target_o, read_target_c_o, sp_mat_index_o,  n_o, k_o, m_o, mem_busy_o);



	// PARAMERES
    parameter DATA_WIDTH = 16; // width of the data BUS in bits
	parameter BUS_WIDTH = 64; // width of the BUS in bits
	parameter ADDR_WIDTH = 16; // width of addres BUS in bits
	localparam MAX_DIM = BUS_WIDTH/DATA_WIDTH; // max dimension of the matrix
	parameter SP_NTARGETS = 4; // number of optionally matrix targets in ScratchPad 
	
	input wire clk_i; // clock
	input wire rst_ni; // reset

	input wire [ADDR_WIDTH-1:0] addr_i; // 
	input wire [BUS_WIDTH-1:0] wdata_i;
	input wire write_i; // write signal from the apb module
	input wire read_i; // read signal from the apb module

	input wire [BUS_WIDTH-1:0] sp_mat_i; // matrix element that arrives from ScratchPad module
	input wire [MAX_DIM**2-1:0] flags_adder_i; // vector of carries that arrives from the Adder module
	input wire [MAX_DIM**2-1:0] flags_systolic_i; // vector of carries that arrives from the systolic array module
	input wire write_flag_i; // signal from the control that tells to write the carries to the flags register
	input wire [MAX_DIM-1:0] strb_i;


	output reg [BUS_WIDTH-1:0] rdata_o; // transfer element from this module to the APB module
	output wire mod_o; // tells the Adder module which operation to execute
	
	output wire [BUS_WIDTH*MAX_DIM-1:0] operand_A_o; // the first operand to multiply - assigned to the buffers module
	output wire [BUS_WIDTH*MAX_DIM-1:0] operand_B_o; // the second operand to multiply - assigned to the buffers module
	
	output reg [SP_NTARGETS/4:0] sp_read_target_o; // the target to read from ScratchPad
	output reg sp_read_o; // read from the ScratchPad
	output wire [MAX_DIM-1:0] sp_mat_index_o;
	
	output wire start_FMEM_o; // tells the control to start the multiply operation
	output wire [1:0] write_target_o; // tells the control what is the target to write in ScratchPad
	output wire [1:0] read_target_c_o; // tells the control what is the target to read from the ScratchPad as Matrix C

	output wire [1:0] n_o;
	output wire [1:0] k_o;
	output wire [1:0] m_o;
	
	output wire mem_busy_o;
	
	reg [15:0] control; // control register
	reg [DATA_WIDTH*MAX_DIM-1:0] matA [MAX_DIM-1:0]; // register that contains Matrix A
	reg [DATA_WIDTH*MAX_DIM-1:0] matB [MAX_DIM-1:0]; // register that contains Matrix B
	reg [MAX_DIM**2-1:0] flags; // register that contains the union of the carries vectors(from systolic array and Adder modules)
	reg rststart;
	reg [3:0] busy_line;

	wire [MAX_DIM/4:0] mat_index; // index to operate(read/write) in Matrix
	
	integer i;
	integer m; 
	always @(posedge clk_i or negedge rst_ni) begin: CONT
		if(!rst_ni)
		begin
			control <= 0; // clear control register
			for (i=0; i<MAX_DIM; i=i+1) matA[i] <= 0; // clear Matrix A
			for (i=0; i<MAX_DIM; i=i+1) matB[i] <= 0; // clear Matrix B
			flags <= 0; // clear register of carries
			rststart <= 0;
			busy_line <= 0;
		end
		else
		begin
			
			rststart <= control[0];
      
			if((write_i && addr_i[4:0] == 5'b00000) || rststart == 1) // conditions to write to the local registers
			begin
				if(rststart == 1)
					control[0] <= 0;
				else
					control[0] <= wdata_i[0];
				control[15:1] <= wdata_i[15:1]; // write from the apb module to the control register
			end
			if(write_i && addr_i[4:0] == 5'b00100) // conditions to write to the local registers
			begin
			  for(m=0;m<MAX_DIM;m=m+1)
			  begin
			    if(strb_i[m] == 1'b1)
				    matA[mat_index][DATA_WIDTH*(m+1)-1 -:DATA_WIDTH] <= wdata_i[DATA_WIDTH*(m+1)-1 -:DATA_WIDTH]; // write from the apb module to the Matrix A register
				end
			end
			if(write_i && addr_i[4:0] == 5'b01000) // conditions to write to the local registers
			begin
				for(m=0;m<MAX_DIM;m=m+1)
			  begin
			    if(strb_i[m] == 1'b1)
				    matB[mat_index][DATA_WIDTH*(m+1)-1 -:DATA_WIDTH] <= wdata_i[DATA_WIDTH*(m+1)-1 -:DATA_WIDTH]; // write from the apb module to the Matrix B register
				end
			end
			if(write_flag_i) // conditions to write to the local registers
			begin
				flags <= flags_adder_i | flags_systolic_i; // final carries register is generated by the OR operation between 2 carries vectors 
			end
			
			if (write_i && addr_i[4:0] == 5'b00000 && wdata_i[0] == 1)
			begin
			  busy_line <= 4'b1111;
			end
			else
			begin
			  busy_line[3] <= 0;
			  busy_line[2] <= busy_line[3];
			  busy_line[1] <= busy_line[2];
			  busy_line[0] <= busy_line[1];
			end
		end
	end
	
	always @*
	begin:RDATA_ASSIGN
	  rdata_o = 0;
		if(read_i) // read request from the apb module
		begin
		
			case(addr_i[4:0]) // export data to apb via address 
			5'b00000: 
				rdata_o = {{(BUS_WIDTH-16){1'b0}}, control}; // export control register to apb module
			5'b00100:
				rdata_o = matA[mat_index]; // export element of Matrix A to the apb module
			5'b01000:
				rdata_o = matB[mat_index]; // export element of Matrix B to the apb module
			5'b01100:
				rdata_o = {{(BUS_WIDTH-MAX_DIM**2){1'b0}}, flags}; // export the carries register to the apb module
			5'b10000:
				rdata_o = sp_mat_i; // export dedicated element of chosen matrix from ScratchPad module 
			5'b10100:
				rdata_o = sp_mat_i; // export dedicated element of chosen matrix from ScratchPad module 
			5'b11000:
				rdata_o = sp_mat_i; // export dedicated element of chosen matrix from ScratchPad module 
			5'b11100:
				rdata_o = sp_mat_i; // export dedicated element of chosen matrix from ScratchPad module 
			default:
				rdata_o = 0;
			endcase
		end
	end


	case(SP_NTARGETS)
	// case of 4 matrixes targets in ScratchPad
	4: begin
		always @*
		begin: sp_addr
			case(addr_i[4:0])
			5'b10000:
				sp_read_target_o = 2'b00; // first target to read from the ScratchPad
			5'b10100:
				sp_read_target_o = 2'b01; // second target to read from the ScratchPad
			5'b11000:
				sp_read_target_o = 2'b10; // third target to read from the ScratchPad
			5'b11100:
				sp_read_target_o = 2'b11; // fourth target to read from the ScratchPad
			default:
				sp_read_target_o = 2'b00;
			endcase
			
		end
	end
	// case of 2 matrixes targets in ScratchPad
	2: begin
		always @*
		begin: sp_addr
			case(addr_i[4:0])
			5'b10000:
				sp_read_target_o = 1'b0; // first target to read from the ScratchPad
			5'b10100:
				sp_read_target_o = 1'b1; // second target to read from the ScratchPad
			default:
				sp_read_target_o = 1'b0;
			endcase
			
		end
	end
	// case of 1 matrixes target in ScratchPad
	1: begin
		always @*
		begin: sp_addr
			sp_read_target_o = 1'b0; // target to read from the ScratchPad
		end
		end
	endcase



	case(SP_NTARGETS)
	// case of 4 matrixes targets in ScratchPad
	4: begin
		always @*
		begin: sp_reado
			if(read_i && (addr_i[4:0] == 5'b10000 || addr_i[4:0] == 5'b10100 || addr_i[4:0] == 5'b11000 || addr_i[4:0] == 5'b11100)) // conditions to read to the local registers from the ScratchPad module
				sp_read_o = 1'b1;
			else
				sp_read_o = 1'b0;
		end
	end
	// case of 2 matrixes targets in ScratchPad
	2: begin
		always @*
		begin: sp_reado
			if(read_i && (addr_i[4:0] == 5'b10000 || addr_i[4:0] == 5'b10100)) // conditions to read to the local registers from the ScratchPad module
				sp_read_o = 1'b1;
			else
				sp_read_o = 1'b0;
		end
	end
	// case of 1 matrix targets in ScratchPad
	1: begin
		always @*
		begin: sp_reado
			if(read_i && addr_i[4:0] == 5'b10000) // conditions to read to the local registers from the ScratchPad module
				sp_read_o = 1'b1;
			else
				sp_read_o = 1'b0;
		end
		end
	endcase


	generate
	case(MAX_DIM)
	4: assign mat_index = addr_i[6:5]; // sub - addressing (in case of 4 we need 2 bit)
	default: assign mat_index = addr_i[5]; // sub - addressing (in case of 1,2 we need 1 bit)
	endcase
	endgenerate

	generate
	case(MAX_DIM)
	4: assign sp_mat_index_o = addr_i[8:5];//ביטים בעיה
	2: assign sp_mat_index_o = addr_i[6:5]; // sub - addressing (in case of 4 we need 2 bit)
	default: assign sp_mat_index_o = addr_i[5]; // sub - addressing (in case of 1,2 we need 1 bit)
	endcase
	endgenerate


	assign start_FMEM_o = control[0]; // start bit - connected to the control module
	assign mod_o = control[1]; // mod bit - connected to the control and Adder modules
	assign write_target_o = control[3:2]; // matrix write target - connected to the control (the final target is in the ScratchPad)
	assign read_target_c_o = control[5:4];// matrix C read target - connected to the control (the final target is in the ScratchPad)
	assign n_o = control[9:8];
	assign k_o = control[11:10];
	assign m_o = control[13:12];
	assign mem_busy_o = busy_line[0];

	genvar j;
	generate
	for (j=0; j<MAX_DIM; j=j+1)
		assign operand_A_o[BUS_WIDTH*(j+1)-1 -:BUS_WIDTH] = matA[j]; // assisn the register of matrix A to the output => buffers nodule
	endgenerate
	generate
	for (j=0; j<MAX_DIM; j=j+1)
		assign operand_B_o[BUS_WIDTH*(j+1)-1 -:BUS_WIDTH] = matB[j]; // assisn the register of matrix B to the output => buffers nodule
	endgenerate

endmodule
